module line(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h0c000006;
30'h00000002: inst = 32'h37bd4000;
30'h00000003: inst = 32'h3c0c4000;
30'h00000004: inst = 32'h01800008;
30'h00000005: inst = 32'h00000000;
30'h00000006: inst = 32'h27bdffe8;
30'h00000007: inst = 32'h3c021900;
30'h00000008: inst = 32'h3c030100;
30'h00000009: inst = 32'h3c0402ff;
30'h0000000a: inst = 32'h34450000;
30'h0000000b: inst = 32'h34660000;
30'h0000000c: inst = 32'hafa00010;
30'h0000000d: inst = 32'h3487ff0f;
30'h0000000e: inst = 32'h34480004;
30'h0000000f: inst = 32'haca60000;
30'h00000010: inst = 32'h3c090320;
30'h00000011: inst = 32'h240a0060;
30'h00000012: inst = 32'h344b0008;
30'h00000013: inst = 32'had070000;
30'h00000014: inst = 32'h3c070200;
30'h00000015: inst = 32'h35280060;
30'h00000016: inst = 32'h344c000c;
30'h00000017: inst = 32'had6a0000;
30'h00000018: inst = 32'h34eaffff;
30'h00000019: inst = 32'h344b0010;
30'h0000001a: inst = 32'had880000;
30'h0000001b: inst = 32'h24080200;
30'h0000001c: inst = 32'h344c0014;
30'h0000001d: inst = 32'had6a0000;
30'h0000001e: inst = 32'h352a0200;
30'h0000001f: inst = 32'h344b0018;
30'h00000020: inst = 32'had880000;
30'h00000021: inst = 32'h34e800ff;
30'h00000022: inst = 32'h344c001c;
30'h00000023: inst = 32'had6a0000;
30'h00000024: inst = 32'h240a012c;
30'h00000025: inst = 32'h344b0020;
30'h00000026: inst = 32'had880000;
30'h00000027: inst = 32'h3528012c;
30'h00000028: inst = 32'h344c0024;
30'h00000029: inst = 32'had6a0000;
30'h0000002a: inst = 32'h348a00ff;
30'h0000002b: inst = 32'h344b0028;
30'h0000002c: inst = 32'had880000;
30'h0000002d: inst = 32'h24080100;
30'h0000002e: inst = 32'h344c002c;
30'h0000002f: inst = 32'had6a0000;
30'h00000030: inst = 32'h352a0100;
30'h00000031: inst = 32'h344b0030;
30'h00000032: inst = 32'had880000;
30'h00000033: inst = 32'h3c0801a0;
30'h00000034: inst = 32'h348cff00;
30'h00000035: inst = 32'h344d0034;
30'h00000036: inst = 32'had6a0000;
30'h00000037: inst = 32'h350a0000;
30'h00000038: inst = 32'h344b0038;
30'h00000039: inst = 32'hadac0000;
30'h0000003a: inst = 32'h35080258;
30'h0000003b: inst = 32'h344c003c;
30'h0000003c: inst = 32'had6a0000;
30'h0000003d: inst = 32'h3c0a01b0;
30'h0000003e: inst = 32'h348b0000;
30'h0000003f: inst = 32'h344d0040;
30'h00000040: inst = 32'had880000;
30'h00000041: inst = 32'h35480000;
30'h00000042: inst = 32'h344c0044;
30'h00000043: inst = 32'hadab0000;
30'h00000044: inst = 32'h354a0258;
30'h00000045: inst = 32'h344b0048;
30'h00000046: inst = 32'had880000;
30'h00000047: inst = 32'h34e7ff00;
30'h00000048: inst = 32'h3448004c;
30'h00000049: inst = 32'had6a0000;
30'h0000004a: inst = 32'h344a0050;
30'h0000004b: inst = 32'had070000;
30'h0000004c: inst = 32'h34630258;
30'h0000004d: inst = 32'h34470054;
30'h0000004e: inst = 32'had460000;
30'h0000004f: inst = 32'h3484ffff;
30'h00000050: inst = 32'h34460058;
30'h00000051: inst = 32'hace30000;
30'h00000052: inst = 32'h3443005c;
30'h00000053: inst = 32'hacc40000;
30'h00000054: inst = 32'h35240000;
30'h00000055: inst = 32'h34460060;
30'h00000056: inst = 32'hac600000;
30'h00000057: inst = 32'h3c031800;
30'h00000058: inst = 32'h3c071040;
30'h00000059: inst = 32'h34420064;
30'h0000005a: inst = 32'hacc40000;
30'h0000005b: inst = 32'h34e40000;
30'h0000005c: inst = 32'h34660004;
30'h0000005d: inst = 32'hac400000;
30'h0000005e: inst = 32'h34620000;
30'h0000005f: inst = 32'hacc40000;
30'h00000060: inst = 32'hac450000;
30'h00000061: inst = 32'h24020000;
30'h00000062: inst = 32'h27bd0018;
30'h00000063: inst = 32'h03e00008;
30'h00000064: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
