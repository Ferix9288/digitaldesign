module demo(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h37bd4000;
30'h00000002: inst = 32'h3c011fff;
30'h00000003: inst = 32'hac20001c;
30'h00000004: inst = 32'h3c011fff;
30'h00000005: inst = 32'hac200020;
30'h00000006: inst = 32'h3c011bef;
30'h00000007: inst = 32'hac28f000;
30'h00000008: inst = 32'h3c011fff;
30'h00000009: inst = 32'hac200028;
30'h0000000a: inst = 32'h24090001;
30'h0000000b: inst = 32'h3c011fff;
30'h0000000c: inst = 32'hac200030;
30'h0000000d: inst = 32'h3c011fff;
30'h0000000e: inst = 32'hac200034;
30'h0000000f: inst = 32'h3c0802fa;
30'h00000010: inst = 32'h3508f000;
30'h00000011: inst = 32'h40884800;
30'h00000012: inst = 32'h3c0902fa;
30'h00000013: inst = 32'h3529f080;
30'h00000014: inst = 32'h40895800;
30'h00000015: inst = 32'h340afc01;
30'h00000016: inst = 32'h408a6000;
30'h00000017: inst = 32'h0c000048;
30'h00000018: inst = 32'h00000000;
30'h00000019: inst = 32'h27bdffe0;
30'h0000001a: inst = 32'hafa40010;
30'h0000001b: inst = 32'hafa50014;
30'h0000001c: inst = 32'hafa60018;
30'h0000001d: inst = 32'h8fa20010;
30'h0000001e: inst = 32'h00000000;
30'h0000001f: inst = 32'h8c430000;
30'h00000020: inst = 32'h00000000;
30'h00000021: inst = 32'h8fa40014;
30'h00000022: inst = 32'h00000000;
30'h00000023: inst = 32'h00641821;
30'h00000024: inst = 32'hac430000;
30'h00000025: inst = 32'h8fa20010;
30'h00000026: inst = 32'h00000000;
30'h00000027: inst = 32'h8c430004;
30'h00000028: inst = 32'h00000000;
30'h00000029: inst = 32'h8fa40018;
30'h0000002a: inst = 32'h00000000;
30'h0000002b: inst = 32'h3c051780;
30'h0000002c: inst = 32'h3c060100;
30'h0000002d: inst = 32'h00641821;
30'h0000002e: inst = 32'h3c0403ff;
30'h0000002f: inst = 32'h34c60000;
30'h00000030: inst = 32'h34a70000;
30'h00000031: inst = 32'hac430004;
30'h00000032: inst = 32'h3482ffff;
30'h00000033: inst = 32'h34a30004;
30'h00000034: inst = 32'hace60000;
30'h00000035: inst = 32'hac620000;
30'h00000036: inst = 32'h8fa20010;
30'h00000037: inst = 32'h00000000;
30'h00000038: inst = 32'h8c430004;
30'h00000039: inst = 32'h00000000;
30'h0000003a: inst = 32'h8c420000;
30'h0000003b: inst = 32'h00000000;
30'h0000003c: inst = 32'h00031b00;
30'h0000003d: inst = 32'h00021580;
30'h0000003e: inst = 32'h00621021;
30'h0000003f: inst = 32'h3442000a;
30'h00000040: inst = 32'h34a30008;
30'h00000041: inst = 32'h34a4000c;
30'h00000042: inst = 32'hac620000;
30'h00000043: inst = 32'hac800000;
30'h00000044: inst = 32'h24020000;
30'h00000045: inst = 32'h27bd0020;
30'h00000046: inst = 32'h03e00008;
30'h00000047: inst = 32'h00000000;
30'h00000048: inst = 32'h27bdffb8;
30'h00000049: inst = 32'hafbf0044;
30'h0000004a: inst = 32'h3c021000;
30'h0000004b: inst = 32'h244202b0;
30'h0000004c: inst = 32'hafa00020;
30'h0000004d: inst = 32'h8c430000;
30'h0000004e: inst = 32'h00000000;
30'h0000004f: inst = 32'h8c420004;
30'h00000050: inst = 32'h00000000;
30'h00000051: inst = 32'hafa30038;
30'h00000052: inst = 32'hafa2003c;
30'h00000053: inst = 32'h3c021bee;
30'h00000054: inst = 32'h24030001;
30'h00000055: inst = 32'h3442f000;
30'h00000056: inst = 32'hafa30034;
30'h00000057: inst = 32'h8c420000;
30'h00000058: inst = 32'h00000000;
30'h00000059: inst = 32'h24030072;
30'h0000005a: inst = 32'h0062182a;
30'h0000005b: inst = 32'h1460000b;
30'h0000005c: inst = 32'h00000000;
30'h0000005d: inst = 32'h24030061;
30'h0000005e: inst = 32'h10430015;
30'h0000005f: inst = 32'h00000000;
30'h00000060: inst = 32'h24030064;
30'h00000061: inst = 32'h14430020;
30'h00000062: inst = 32'h00000000;
30'h00000063: inst = 32'h27a40038;
30'h00000064: inst = 32'h24050001;
30'h00000065: inst = 32'h08000076;
30'h00000066: inst = 32'h00000000;
30'h00000067: inst = 32'h24030073;
30'h00000068: inst = 32'h10430012;
30'h00000069: inst = 32'h00000000;
30'h0000006a: inst = 32'h24030077;
30'h0000006b: inst = 32'h14430016;
30'h0000006c: inst = 32'h00000000;
30'h0000006d: inst = 32'h27a40038;
30'h0000006e: inst = 32'h24050000;
30'h0000006f: inst = 32'h2406ffff;
30'h00000070: inst = 32'h0c000019;
30'h00000071: inst = 32'h00000000;
30'h00000072: inst = 32'h08000083;
30'h00000073: inst = 32'h00000000;
30'h00000074: inst = 32'h27a40038;
30'h00000075: inst = 32'h2405ffff;
30'h00000076: inst = 32'h24060000;
30'h00000077: inst = 32'h0c000019;
30'h00000078: inst = 32'h00000000;
30'h00000079: inst = 32'h08000083;
30'h0000007a: inst = 32'h00000000;
30'h0000007b: inst = 32'h27a40038;
30'h0000007c: inst = 32'h24050000;
30'h0000007d: inst = 32'h24060001;
30'h0000007e: inst = 32'h0c000019;
30'h0000007f: inst = 32'h00000000;
30'h00000080: inst = 32'h08000083;
30'h00000081: inst = 32'h00000000;
30'h00000082: inst = 32'hafa00034;
30'h00000083: inst = 32'h8fa20034;
30'h00000084: inst = 32'h00000000;
30'h00000085: inst = 32'h10400016;
30'h00000086: inst = 32'h00000000;
30'h00000087: inst = 32'h3c020800;
30'h00000088: inst = 32'h34420020;
30'h00000089: inst = 32'h3c031040;
30'h0000008a: inst = 32'h8c420000;
30'h0000008b: inst = 32'h00000000;
30'h0000008c: inst = 32'h34630000;
30'h0000008d: inst = 32'h14430004;
30'h0000008e: inst = 32'h00000000;
30'h0000008f: inst = 32'h3c021080;
30'h00000090: inst = 32'h08000093;
30'h00000091: inst = 32'h00000000;
30'h00000092: inst = 32'h3c021040;
30'h00000093: inst = 32'h3c031800;
30'h00000094: inst = 32'h34420000;
30'h00000095: inst = 32'h34630004;
30'h00000096: inst = 32'hac620000;
30'h00000097: inst = 32'h3c028000;
30'h00000098: inst = 32'h8fa30028;
30'h00000099: inst = 32'h00000000;
30'h0000009a: inst = 32'h34420040;
30'h0000009b: inst = 32'hac430000;
30'h0000009c: inst = 32'h3c020800;
30'h0000009d: inst = 32'h34420020;
30'h0000009e: inst = 32'h8c420000;
30'h0000009f: inst = 32'h00000000;
30'h000000a0: inst = 32'hafa20030;
30'h000000a1: inst = 32'h3c020800;
30'h000000a2: inst = 32'h34420020;
30'h000000a3: inst = 32'h8c420000;
30'h000000a4: inst = 32'h00000000;
30'h000000a5: inst = 32'h8fa30030;
30'h000000a6: inst = 32'h00000000;
30'h000000a7: inst = 32'h1043fff9;
30'h000000a8: inst = 32'h00000000;
30'h000000a9: inst = 32'h08000053;
30'h000000aa: inst = 32'h00000000;
30'h000000ab: inst = 32'h00000000;
30'h000000ac: inst = 32'h00000190;
30'h000000ad: inst = 32'h00000226;
default:      inst = 32'h00000000;
endcase
end
endmodule
