module fifo(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d0100;
30'h00000001: inst = 32'h0ffffc79;
30'h00000002: inst = 32'h37bd3000;
30'h00000003: inst = 32'h27bdffe8;
30'h00000004: inst = 32'h3c028000;
30'h00000005: inst = 32'hafa40010;
30'h00000006: inst = 32'h34420000;
30'h00000007: inst = 32'hafa00014;
30'h00000008: inst = 32'h8c420000;
30'h00000009: inst = 32'h00000000;
30'h0000000a: inst = 32'h30420001;
30'h0000000b: inst = 32'h1040000b;
30'h0000000c: inst = 32'h00000000;
30'h0000000d: inst = 32'h8fa20014;
30'h0000000e: inst = 32'h00000000;
30'h0000000f: inst = 32'h8fa30010;
30'h00000010: inst = 32'h00000000;
30'h00000011: inst = 32'h00621021;
30'h00000012: inst = 32'h80420000;
30'h00000013: inst = 32'h00000000;
30'h00000014: inst = 32'h3c038000;
30'h00000015: inst = 32'h34630008;
30'h00000016: inst = 32'hac620000;
30'h00000017: inst = 32'h8fa20014;
30'h00000018: inst = 32'h00000000;
30'h00000019: inst = 32'h8fa30010;
30'h0000001a: inst = 32'h00000000;
30'h0000001b: inst = 32'h00621021;
30'h0000001c: inst = 32'h3c031fff;
30'h0000001d: inst = 32'h90420000;
30'h0000001e: inst = 32'h00000000;
30'h0000001f: inst = 32'h34640015;
30'h00000020: inst = 32'h34630000;
30'h00000021: inst = 32'h8c840000;
30'h00000022: inst = 32'h00000000;
30'h00000023: inst = 32'h00831821;
30'h00000024: inst = 32'ha0620000;
30'h00000025: inst = 32'h90620000;
30'h00000026: inst = 32'h00000000;
30'h00000027: inst = 32'h14400004;
30'h00000028: inst = 32'h00000000;
30'h00000029: inst = 32'h24020000;
30'h0000002a: inst = 32'h0bfffc36;
30'h0000002b: inst = 32'h00000000;
30'h0000002c: inst = 32'h3c021fff;
30'h0000002d: inst = 32'h34430015;
30'h0000002e: inst = 32'h34420016;
30'h0000002f: inst = 32'h8c630000;
30'h00000030: inst = 32'h00000000;
30'h00000031: inst = 32'h8c420000;
30'h00000032: inst = 32'h00000000;
30'h00000033: inst = 32'h2442ffff;
30'h00000034: inst = 32'h00621026;
30'h00000035: inst = 32'h0002102b;
30'h00000036: inst = 32'h30420001;
30'h00000037: inst = 32'h10400016;
30'h00000038: inst = 32'h00000000;
30'h00000039: inst = 32'h3c021fff;
30'h0000003a: inst = 32'h34420015;
30'h0000003b: inst = 32'h3c03cccc;
30'h0000003c: inst = 32'h8c440000;
30'h0000003d: inst = 32'h00000000;
30'h0000003e: inst = 32'h24840001;
30'h0000003f: inst = 32'h3463cccd;
30'h00000040: inst = 32'h00830019;
30'h00000041: inst = 32'h00001810;
30'h00000042: inst = 32'h00031902;
30'h00000043: inst = 32'h24050014;
30'h00000044: inst = 32'h00650018;
30'h00000045: inst = 32'h00001812;
30'h00000046: inst = 32'h00831823;
30'h00000047: inst = 32'hac430000;
30'h00000048: inst = 32'h8fa20014;
30'h00000049: inst = 32'h00000000;
30'h0000004a: inst = 32'h24420001;
30'h0000004b: inst = 32'hafa20014;
30'h0000004c: inst = 32'h0bfffc17;
30'h0000004d: inst = 32'h00000000;
30'h0000004e: inst = 32'h27bd0018;
30'h0000004f: inst = 32'h03e00008;
30'h00000050: inst = 32'h00000000;
30'h00000051: inst = 32'h27bdffe8;
30'h00000052: inst = 32'h3c021fff;
30'h00000053: inst = 32'h34430015;
30'h00000054: inst = 32'h8c630000;
30'h00000055: inst = 32'h00000000;
30'h00000056: inst = 32'h34420016;
30'h00000057: inst = 32'h8c420000;
30'h00000058: inst = 32'h00000000;
30'h00000059: inst = 32'h1062001c;
30'h0000005a: inst = 32'h00000000;
30'h0000005b: inst = 32'h3c021fff;
30'h0000005c: inst = 32'h34430016;
30'h0000005d: inst = 32'h34420000;
30'h0000005e: inst = 32'h8c640000;
30'h0000005f: inst = 32'h00000000;
30'h00000060: inst = 32'h00821021;
30'h00000061: inst = 32'h90420000;
30'h00000062: inst = 32'h00000000;
30'h00000063: inst = 32'ha3a20010;
30'h00000064: inst = 32'h3c028000;
30'h00000065: inst = 32'h83a40010;
30'h00000066: inst = 32'h00000000;
30'h00000067: inst = 32'h34420008;
30'h00000068: inst = 32'hac440000;
30'h00000069: inst = 32'h3c02cccc;
30'h0000006a: inst = 32'h8c640000;
30'h0000006b: inst = 32'h00000000;
30'h0000006c: inst = 32'h24840001;
30'h0000006d: inst = 32'h3442cccd;
30'h0000006e: inst = 32'h00820019;
30'h0000006f: inst = 32'h00001010;
30'h00000070: inst = 32'h00021102;
30'h00000071: inst = 32'h24050014;
30'h00000072: inst = 32'h00450018;
30'h00000073: inst = 32'h00001012;
30'h00000074: inst = 32'h00821023;
30'h00000075: inst = 32'hac620000;
30'h00000076: inst = 32'h27bd0018;
30'h00000077: inst = 32'h03e00008;
30'h00000078: inst = 32'h00000000;
30'h00000079: inst = 32'h27bdffe8;
30'h0000007a: inst = 32'hafa00010;
30'h0000007b: inst = 32'h24020000;
30'h0000007c: inst = 32'h27bd0018;
30'h0000007d: inst = 32'h03e00008;
30'h0000007e: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
