module line(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h0c000006;
30'h00000002: inst = 32'h37bd4000;
30'h00000003: inst = 32'h3c0c4000;
30'h00000004: inst = 32'h01800008;
30'h00000005: inst = 32'h00000000;
30'h00000006: inst = 32'h27bdffe8;
30'h00000007: inst = 32'h3c021900;
30'h00000008: inst = 32'h3c030100;
30'h00000009: inst = 32'h3c040200;
30'h0000000a: inst = 32'h34450000;
30'h0000000b: inst = 32'h34630000;
30'h0000000c: inst = 32'hafa00010;
30'h0000000d: inst = 32'h348600ff;
30'h0000000e: inst = 32'h34470004;
30'h0000000f: inst = 32'haca30000;
30'h00000010: inst = 32'h3c030320;
30'h00000011: inst = 32'h24080258;
30'h00000012: inst = 32'h34490008;
30'h00000013: inst = 32'hace60000;
30'h00000014: inst = 32'h3c0602ff;
30'h00000015: inst = 32'h34670000;
30'h00000016: inst = 32'h344a000c;
30'h00000017: inst = 32'had280000;
30'h00000018: inst = 32'h34c80000;
30'h00000019: inst = 32'h34490010;
30'h0000001a: inst = 32'had470000;
30'h0000001b: inst = 32'h2407012c;
30'h0000001c: inst = 32'h344a0014;
30'h0000001d: inst = 32'had280000;
30'h0000001e: inst = 32'h3468012c;
30'h0000001f: inst = 32'h34490018;
30'h00000020: inst = 32'had470000;
30'h00000021: inst = 32'h3484ff00;
30'h00000022: inst = 32'h34470028;
30'h00000023: inst = 32'had280000;
30'h00000024: inst = 32'h3448002c;
30'h00000025: inst = 32'hace40000;
30'h00000026: inst = 32'h34630258;
30'h00000027: inst = 32'h34440030;
30'h00000028: inst = 32'had000000;
30'h00000029: inst = 32'h3c070190;
30'h0000002a: inst = 32'h34c6ffff;
30'h0000002b: inst = 32'h3448001c;
30'h0000002c: inst = 32'hac830000;
30'h0000002d: inst = 32'h34e30000;
30'h0000002e: inst = 32'h34440020;
30'h0000002f: inst = 32'had060000;
30'h00000030: inst = 32'h34e60258;
30'h00000031: inst = 32'h34470024;
30'h00000032: inst = 32'hac830000;
30'h00000033: inst = 32'h3c031800;
30'h00000034: inst = 32'h3c041040;
30'h00000035: inst = 32'h34420034;
30'h00000036: inst = 32'hace60000;
30'h00000037: inst = 32'h34840000;
30'h00000038: inst = 32'h34660004;
30'h00000039: inst = 32'hac400000;
30'h0000003a: inst = 32'h34620000;
30'h0000003b: inst = 32'hacc40000;
30'h0000003c: inst = 32'hac450000;
30'h0000003d: inst = 32'h24020000;
30'h0000003e: inst = 32'h27bd0018;
30'h0000003f: inst = 32'h03e00008;
30'h00000040: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
