module demo(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h0c000057;
30'h00000002: inst = 32'h37bd4000;
30'h00000003: inst = 32'h27bdffe8;
30'h00000004: inst = 32'h3c021800;
30'h00000005: inst = 32'h34420008;
30'h00000006: inst = 32'h8c430000;
30'h00000007: inst = 32'h00000000;
30'h00000008: inst = 32'h3c041780;
30'h00000009: inst = 32'h3c050200;
30'h0000000a: inst = 32'h24630001;
30'h0000000b: inst = 32'h34a500ff;
30'h0000000c: inst = 32'h34860004;
30'h0000000d: inst = 32'hac430000;
30'h0000000e: inst = 32'hacc50000;
30'h0000000f: inst = 32'h8c430000;
30'h00000010: inst = 32'h00000000;
30'h00000011: inst = 32'h24630020;
30'h00000012: inst = 32'h3c05001a;
30'h00000013: inst = 32'h00031c00;
30'h00000014: inst = 32'h34860008;
30'h00000015: inst = 32'h3c0702ff;
30'h00000016: inst = 32'h34a5002b;
30'h00000017: inst = 32'h3488000c;
30'h00000018: inst = 32'hacc30000;
30'h00000019: inst = 32'h3c031230;
30'h0000001a: inst = 32'h34e60000;
30'h0000001b: inst = 32'h34870010;
30'h0000001c: inst = 32'had050000;
30'h0000001d: inst = 32'h34631234;
30'h0000001e: inst = 32'h34850014;
30'h0000001f: inst = 32'hace60000;
30'h00000020: inst = 32'haca30000;
30'h00000021: inst = 32'h8c420000;
30'h00000022: inst = 32'h00000000;
30'h00000023: inst = 32'h244200aa;
30'h00000024: inst = 32'h34830018;
30'h00000025: inst = 32'h3484001c;
30'h00000026: inst = 32'hac620000;
30'h00000027: inst = 32'hac800000;
30'h00000028: inst = 32'h8fa20010;
30'h00000029: inst = 32'h00000000;
30'h0000002a: inst = 32'h27bd0018;
30'h0000002b: inst = 32'h03e00008;
30'h0000002c: inst = 32'h00000000;
30'h0000002d: inst = 32'h27bdffe8;
30'h0000002e: inst = 32'h3c021800;
30'h0000002f: inst = 32'h34420008;
30'h00000030: inst = 32'h8c430000;
30'h00000031: inst = 32'h00000000;
30'h00000032: inst = 32'h3c041780;
30'h00000033: inst = 32'h3c050200;
30'h00000034: inst = 32'h24630001;
30'h00000035: inst = 32'h34a500ff;
30'h00000036: inst = 32'h34860004;
30'h00000037: inst = 32'hac430000;
30'h00000038: inst = 32'hacc50000;
30'h00000039: inst = 32'h8c430000;
30'h0000003a: inst = 32'h00000000;
30'h0000003b: inst = 32'h24630020;
30'h0000003c: inst = 32'h3c05001a;
30'h0000003d: inst = 32'h00031c00;
30'h0000003e: inst = 32'h34860008;
30'h0000003f: inst = 32'h3c0702ff;
30'h00000040: inst = 32'h34a5002b;
30'h00000041: inst = 32'h3488000c;
30'h00000042: inst = 32'hacc30000;
30'h00000043: inst = 32'h3c031230;
30'h00000044: inst = 32'h34e60000;
30'h00000045: inst = 32'h34870010;
30'h00000046: inst = 32'had050000;
30'h00000047: inst = 32'h34631234;
30'h00000048: inst = 32'h34850014;
30'h00000049: inst = 32'hace60000;
30'h0000004a: inst = 32'haca30000;
30'h0000004b: inst = 32'h8c420000;
30'h0000004c: inst = 32'h00000000;
30'h0000004d: inst = 32'h244200aa;
30'h0000004e: inst = 32'h34830018;
30'h0000004f: inst = 32'h3484001c;
30'h00000050: inst = 32'hac620000;
30'h00000051: inst = 32'hac800000;
30'h00000052: inst = 32'h8fa20010;
30'h00000053: inst = 32'h00000000;
30'h00000054: inst = 32'h27bd0018;
30'h00000055: inst = 32'h03e00008;
30'h00000056: inst = 32'h00000000;
30'h00000057: inst = 32'h27bdffc0;
30'h00000058: inst = 32'hafbf003c;
30'h00000059: inst = 32'hafb00028;
30'h0000005a: inst = 32'hafb1002c;
30'h0000005b: inst = 32'hafb20030;
30'h0000005c: inst = 32'hafb30034;
30'h0000005d: inst = 32'h3c028000;
30'h0000005e: inst = 32'h3c030100;
30'h0000005f: inst = 32'h3c041780;
30'h00000060: inst = 32'h3442001c;
30'h00000061: inst = 32'hafa00020;
30'h00000062: inst = 32'h3c051760;
30'h00000063: inst = 32'h34630000;
30'h00000064: inst = 32'h34840000;
30'h00000065: inst = 32'hac400000;
30'h00000066: inst = 32'h3c021800;
30'h00000067: inst = 32'h34a50000;
30'h00000068: inst = 32'hac830000;
30'h00000069: inst = 32'h34420008;
30'h0000006a: inst = 32'h24040010;
30'h0000006b: inst = 32'haca30000;
30'h0000006c: inst = 32'h240300bb;
30'h0000006d: inst = 32'hac440000;
30'h0000006e: inst = 32'hac430000;
30'h0000006f: inst = 32'h3c028000;
30'h00000070: inst = 32'h3442001c;
30'h00000071: inst = 32'h8c420000;
30'h00000072: inst = 32'h00000000;
30'h00000073: inst = 32'h30420001;
30'h00000074: inst = 32'h1040000b;
30'h00000075: inst = 32'h00000000;
30'h00000076: inst = 32'h3c021080;
30'h00000077: inst = 32'h3c031800;
30'h00000078: inst = 32'h3c101780;
30'h00000079: inst = 32'h3c118000;
30'h0000007a: inst = 32'h34520000;
30'h0000007b: inst = 32'h34730004;
30'h0000007c: inst = 32'h0c000003;
30'h0000007d: inst = 32'h00000000;
30'h0000007e: inst = 32'h08000088;
30'h0000007f: inst = 32'h00000000;
30'h00000080: inst = 32'h3c021040;
30'h00000081: inst = 32'h3c031800;
30'h00000082: inst = 32'h3c101760;
30'h00000083: inst = 32'h3c118000;
30'h00000084: inst = 32'h34520000;
30'h00000085: inst = 32'h34730004;
30'h00000086: inst = 32'h0c00002d;
30'h00000087: inst = 32'h00000000;
30'h00000088: inst = 32'h36020000;
30'h00000089: inst = 32'h36230040;
30'h0000008a: inst = 32'hae720000;
30'h0000008b: inst = 32'hac620000;
30'h0000008c: inst = 32'h3c028000;
30'h0000008d: inst = 32'h3442001c;
30'h0000008e: inst = 32'h8c420000;
30'h0000008f: inst = 32'h00000000;
30'h00000090: inst = 32'hafa20024;
30'h00000091: inst = 32'h3c028000;
30'h00000092: inst = 32'h3442001c;
30'h00000093: inst = 32'h8c420000;
30'h00000094: inst = 32'h00000000;
30'h00000095: inst = 32'h8fa30024;
30'h00000096: inst = 32'h00000000;
30'h00000097: inst = 32'h1043fff9;
30'h00000098: inst = 32'h00000000;
30'h00000099: inst = 32'h0800006f;
30'h0000009a: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
