`ifndef GPCOMMANDS
`define CPCOMMANDS
// graphics processor macros
`define STOP 8'h00
`define FILL 8'h01
`define LINE 8'h02
`define CIRCLE 8'h03
`define COLOR_IDX 23:0
`define OPCODE_IDX 31:24
`define X_ADDR 25:16
`define Y_ADDR 9:0

`endif
