module demo(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h37bd4000;
30'h00000002: inst = 32'h3c011fff;
30'h00000003: inst = 32'hac20001c;
30'h00000004: inst = 32'h3c011fff;
30'h00000005: inst = 32'hac200020;
30'h00000006: inst = 32'h24080056;
30'h00000007: inst = 32'h3c011bef;
30'h00000008: inst = 32'hac28f000;
30'h00000009: inst = 32'h3c011fff;
30'h0000000a: inst = 32'hac200028;
30'h0000000b: inst = 32'h24090001;
30'h0000000c: inst = 32'h3c011fff;
30'h0000000d: inst = 32'hac200030;
30'h0000000e: inst = 32'h3c011fff;
30'h0000000f: inst = 32'hac200034;
30'h00000010: inst = 32'h3c0802fa;
30'h00000011: inst = 32'h3508f000;
30'h00000012: inst = 32'h40884800;
30'h00000013: inst = 32'h3c0902fa;
30'h00000014: inst = 32'h3529f080;
30'h00000015: inst = 32'h40895800;
30'h00000016: inst = 32'h340afc01;
30'h00000017: inst = 32'h408a6000;
30'h00000018: inst = 32'h0c0000cb;
30'h00000019: inst = 32'h00000000;
30'h0000001a: inst = 32'h240a0000;
30'h0000001b: inst = 32'h408a6000;
30'h0000001c: inst = 32'h3c0c4000;
30'h0000001d: inst = 32'h01800008;
30'h0000001e: inst = 32'h00000000;
30'h0000001f: inst = 32'h27bdfff0;
30'h00000020: inst = 32'h27bd0010;
30'h00000021: inst = 32'h03e00008;
30'h00000022: inst = 32'h00000000;
30'h00000023: inst = 32'h27bdffc8;
30'h00000024: inst = 32'hafa40014;
30'h00000025: inst = 32'hafa50018;
30'h00000026: inst = 32'hafa6001c;
30'h00000027: inst = 32'h8fa20048;
30'h00000028: inst = 32'h00000000;
30'h00000029: inst = 32'hafa70020;
30'h0000002a: inst = 32'h8fa3004c;
30'h0000002b: inst = 32'h00000000;
30'h0000002c: inst = 32'hafa20024;
30'h0000002d: inst = 32'h8fa20050;
30'h0000002e: inst = 32'h00000000;
30'h0000002f: inst = 32'hafa30028;
30'h00000030: inst = 32'hafa2002c;
30'h00000031: inst = 32'h8fa20018;
30'h00000032: inst = 32'h00000000;
30'h00000033: inst = 32'hafa20030;
30'h00000034: inst = 32'h8fa20018;
30'h00000035: inst = 32'h00000000;
30'h00000036: inst = 32'h8fa30028;
30'h00000037: inst = 32'h00000000;
30'h00000038: inst = 32'h00431021;
30'h00000039: inst = 32'h8fa30030;
30'h0000003a: inst = 32'h00000000;
30'h0000003b: inst = 32'h0043102a;
30'h0000003c: inst = 32'h14400036;
30'h0000003d: inst = 32'h00000000;
30'h0000003e: inst = 32'h3c021bee;
30'h0000003f: inst = 32'h8fa30024;
30'h00000040: inst = 32'h00000000;
30'h00000041: inst = 32'h3442f004;
30'h00000042: inst = 32'h8c440000;
30'h00000043: inst = 32'h00000000;
30'h00000044: inst = 32'h00042080;
30'h00000045: inst = 32'h8fa5002c;
30'h00000046: inst = 32'h00000000;
30'h00000047: inst = 32'h24630002;
30'h00000048: inst = 32'h00a42021;
30'h00000049: inst = 32'hac830000;
30'h0000004a: inst = 32'h8fa30014;
30'h0000004b: inst = 32'h00000000;
30'h0000004c: inst = 32'h8fa40018;
30'h0000004d: inst = 32'h00000000;
30'h0000004e: inst = 32'h8fa50030;
30'h0000004f: inst = 32'h00000000;
30'h00000050: inst = 32'h8c460000;
30'h00000051: inst = 32'h00000000;
30'h00000052: inst = 32'h00852021;
30'h00000053: inst = 32'h24840010;
30'h00000054: inst = 32'h00062880;
30'h00000055: inst = 32'h8fa6002c;
30'h00000056: inst = 32'h00000000;
30'h00000057: inst = 32'h00831804;
30'h00000058: inst = 32'h00a62021;
30'h00000059: inst = 32'hac830004;
30'h0000005a: inst = 32'h8fa3001c;
30'h0000005b: inst = 32'h00000000;
30'h0000005c: inst = 32'h8fa40020;
30'h0000005d: inst = 32'h00000000;
30'h0000005e: inst = 32'h8fa50030;
30'h0000005f: inst = 32'h00000000;
30'h00000060: inst = 32'h8c460000;
30'h00000061: inst = 32'h00000000;
30'h00000062: inst = 32'h00852021;
30'h00000063: inst = 32'h24840010;
30'h00000064: inst = 32'h00062880;
30'h00000065: inst = 32'h8fa6002c;
30'h00000066: inst = 32'h00000000;
30'h00000067: inst = 32'h00831804;
30'h00000068: inst = 32'h00a62021;
30'h00000069: inst = 32'hac830008;
30'h0000006a: inst = 32'h8c430000;
30'h0000006b: inst = 32'h00000000;
30'h0000006c: inst = 32'h24630003;
30'h0000006d: inst = 32'hac430000;
30'h0000006e: inst = 32'h8fa20030;
30'h0000006f: inst = 32'h00000000;
30'h00000070: inst = 32'h24420001;
30'h00000071: inst = 32'h08000033;
30'h00000072: inst = 32'h00000000;
30'h00000073: inst = 32'h3c021bee;
30'h00000074: inst = 32'h3442f004;
30'h00000075: inst = 32'h8c430000;
30'h00000076: inst = 32'h00000000;
30'h00000077: inst = 32'h00031880;
30'h00000078: inst = 32'h8fa4002c;
30'h00000079: inst = 32'h00000000;
30'h0000007a: inst = 32'h00831821;
30'h0000007b: inst = 32'hac600000;
30'h0000007c: inst = 32'h8c430000;
30'h0000007d: inst = 32'h00000000;
30'h0000007e: inst = 32'h24630001;
30'h0000007f: inst = 32'hac430000;
30'h00000080: inst = 32'h27bd0038;
30'h00000081: inst = 32'h03e00008;
30'h00000082: inst = 32'h00000000;
30'h00000083: inst = 32'h27bdffe0;
30'h00000084: inst = 32'hafa40010;
30'h00000085: inst = 32'hafa50014;
30'h00000086: inst = 32'hafa60018;
30'h00000087: inst = 32'hafa7001c;
30'h00000088: inst = 32'h8fa20010;
30'h00000089: inst = 32'h00000000;
30'h0000008a: inst = 32'h8c430000;
30'h0000008b: inst = 32'h00000000;
30'h0000008c: inst = 32'h8fa40014;
30'h0000008d: inst = 32'h00000000;
30'h0000008e: inst = 32'h00641821;
30'h0000008f: inst = 32'hac430000;
30'h00000090: inst = 32'h8fa20010;
30'h00000091: inst = 32'h00000000;
30'h00000092: inst = 32'h8c430004;
30'h00000093: inst = 32'h00000000;
30'h00000094: inst = 32'h8fa40018;
30'h00000095: inst = 32'h00000000;
30'h00000096: inst = 32'h3c051bee;
30'h00000097: inst = 32'h00641821;
30'h00000098: inst = 32'h34a4f004;
30'h00000099: inst = 32'hac430004;
30'h0000009a: inst = 32'h8c820000;
30'h0000009b: inst = 32'h00000000;
30'h0000009c: inst = 32'h3c030100;
30'h0000009d: inst = 32'h00021080;
30'h0000009e: inst = 32'h8fa5001c;
30'h0000009f: inst = 32'h00000000;
30'h000000a0: inst = 32'h34630000;
30'h000000a1: inst = 32'h00a21021;
30'h000000a2: inst = 32'hac430000;
30'h000000a3: inst = 32'h8c820000;
30'h000000a4: inst = 32'h00000000;
30'h000000a5: inst = 32'h3c0303ff;
30'h000000a6: inst = 32'h00021080;
30'h000000a7: inst = 32'h8fa5001c;
30'h000000a8: inst = 32'h00000000;
30'h000000a9: inst = 32'h34630000;
30'h000000aa: inst = 32'h00451021;
30'h000000ab: inst = 32'hac430004;
30'h000000ac: inst = 32'h8fa20010;
30'h000000ad: inst = 32'h00000000;
30'h000000ae: inst = 32'h8c430004;
30'h000000af: inst = 32'h00000000;
30'h000000b0: inst = 32'h8c420000;
30'h000000b1: inst = 32'h00000000;
30'h000000b2: inst = 32'h8c850000;
30'h000000b3: inst = 32'h00000000;
30'h000000b4: inst = 32'h00031b00;
30'h000000b5: inst = 32'h00021580;
30'h000000b6: inst = 32'h00621021;
30'h000000b7: inst = 32'h00051880;
30'h000000b8: inst = 32'h8fa5001c;
30'h000000b9: inst = 32'h00000000;
30'h000000ba: inst = 32'h34420030;
30'h000000bb: inst = 32'h00651821;
30'h000000bc: inst = 32'hac620008;
30'h000000bd: inst = 32'h8c820000;
30'h000000be: inst = 32'h00000000;
30'h000000bf: inst = 32'h00021080;
30'h000000c0: inst = 32'h8fa3001c;
30'h000000c1: inst = 32'h00000000;
30'h000000c2: inst = 32'h00431021;
30'h000000c3: inst = 32'hac40000c;
30'h000000c4: inst = 32'h8c820000;
30'h000000c5: inst = 32'h00000000;
30'h000000c6: inst = 32'h24420004;
30'h000000c7: inst = 32'hac820000;
30'h000000c8: inst = 32'h27bd0020;
30'h000000c9: inst = 32'h03e00008;
30'h000000ca: inst = 32'h00000000;
30'h000000cb: inst = 32'h27bdff98;
30'h000000cc: inst = 32'hafbf0064;
30'h000000cd: inst = 32'hafb00058;
30'h000000ce: inst = 32'hafb1005c;
30'h000000cf: inst = 32'h3c021000;
30'h000000d0: inst = 32'h24420660;
30'h000000d1: inst = 32'hafa0002c;
30'h000000d2: inst = 32'h8c430000;
30'h000000d3: inst = 32'h00000000;
30'h000000d4: inst = 32'h8c420004;
30'h000000d5: inst = 32'h00000000;
30'h000000d6: inst = 32'hafa30050;
30'h000000d7: inst = 32'hafa20054;
30'h000000d8: inst = 32'h3c021780;
30'h000000d9: inst = 32'h3c038000;
30'h000000da: inst = 32'h27a40050;
30'h000000db: inst = 32'h24050000;
30'h000000dc: inst = 32'h34470000;
30'h000000dd: inst = 32'h3c101040;
30'h000000de: inst = 32'h34710020;
30'h000000df: inst = 32'h00053021;
30'h000000e0: inst = 32'h0c000083;
30'h000000e1: inst = 32'h00000000;
30'h000000e2: inst = 32'h36020000;
30'h000000e3: inst = 32'h8e230000;
30'h000000e4: inst = 32'h00000000;
30'h000000e5: inst = 32'h00621826;
30'h000000e6: inst = 32'h3c041080;
30'h000000e7: inst = 32'h2c630001;
30'h000000e8: inst = 32'h34840000;
30'h000000e9: inst = 32'h14600002;
30'h000000ea: inst = 32'h00000000;
30'h000000eb: inst = 32'h00022021;
30'h000000ec: inst = 32'hafa40040;
30'h000000ed: inst = 32'h14820004;
30'h000000ee: inst = 32'h00000000;
30'h000000ef: inst = 32'h3c021780;
30'h000000f0: inst = 32'h080000f3;
30'h000000f1: inst = 32'h00000000;
30'h000000f2: inst = 32'h3c021900;
30'h000000f3: inst = 32'h34420000;
30'h000000f4: inst = 32'h3c031040;
30'h000000f5: inst = 32'hafa20048;
30'h000000f6: inst = 32'h34620000;
30'h000000f7: inst = 32'h8fa30040;
30'h000000f8: inst = 32'h00000000;
30'h000000f9: inst = 32'h00621026;
30'h000000fa: inst = 32'h3c031780;
30'h000000fb: inst = 32'h3c041900;
30'h000000fc: inst = 32'h2c420001;
30'h000000fd: inst = 32'h34630000;
30'h000000fe: inst = 32'h14400002;
30'h000000ff: inst = 32'h00000000;
30'h00000100: inst = 32'h34830000;
30'h00000101: inst = 32'h3c021800;
30'h00000102: inst = 32'hafa30034;
30'h00000103: inst = 32'h8fa30040;
30'h00000104: inst = 32'h00000000;
30'h00000105: inst = 32'h34440004;
30'h00000106: inst = 32'hac830000;
30'h00000107: inst = 32'h3c031bee;
30'h00000108: inst = 32'h8fa40034;
30'h00000109: inst = 32'h00000000;
30'h0000010a: inst = 32'h34420000;
30'h0000010b: inst = 32'h3463f004;
30'h0000010c: inst = 32'hac440000;
30'h0000010d: inst = 32'hac600000;
30'h0000010e: inst = 32'h3c021bee;
30'h0000010f: inst = 32'h3442f004;
30'h00000110: inst = 32'h3c038000;
30'h00000111: inst = 32'h24040001;
30'h00000112: inst = 32'hac400000;
30'h00000113: inst = 32'h3c021040;
30'h00000114: inst = 32'h34630020;
30'h00000115: inst = 32'hafa40044;
30'h00000116: inst = 32'h34420000;
30'h00000117: inst = 32'h8c630000;
30'h00000118: inst = 32'h00000000;
30'h00000119: inst = 32'h00621826;
30'h0000011a: inst = 32'h3c041080;
30'h0000011b: inst = 32'h2c630001;
30'h0000011c: inst = 32'h34840000;
30'h0000011d: inst = 32'h14600002;
30'h0000011e: inst = 32'h00000000;
30'h0000011f: inst = 32'h00022021;
30'h00000120: inst = 32'hafa40040;
30'h00000121: inst = 32'h14820004;
30'h00000122: inst = 32'h00000000;
30'h00000123: inst = 32'h3c021780;
30'h00000124: inst = 32'h08000127;
30'h00000125: inst = 32'h00000000;
30'h00000126: inst = 32'h3c021900;
30'h00000127: inst = 32'h34420000;
30'h00000128: inst = 32'h3c031040;
30'h00000129: inst = 32'hafa20048;
30'h0000012a: inst = 32'h34620000;
30'h0000012b: inst = 32'h8fa30040;
30'h0000012c: inst = 32'h00000000;
30'h0000012d: inst = 32'h00621026;
30'h0000012e: inst = 32'h3c031780;
30'h0000012f: inst = 32'h3c041900;
30'h00000130: inst = 32'h2c420001;
30'h00000131: inst = 32'h34630000;
30'h00000132: inst = 32'h14400002;
30'h00000133: inst = 32'h00000000;
30'h00000134: inst = 32'h34830000;
30'h00000135: inst = 32'hafa30034;
30'h00000136: inst = 32'h3c0200ff;
30'h00000137: inst = 32'h8fa30048;
30'h00000138: inst = 32'h00000000;
30'h00000139: inst = 32'h3442ffff;
30'h0000013a: inst = 32'h24040014;
30'h0000013b: inst = 32'hafa20010;
30'h0000013c: inst = 32'hafa40014;
30'h0000013d: inst = 32'hafa30018;
30'h0000013e: inst = 32'h3c101bee;
30'h0000013f: inst = 32'h24060320;
30'h00000140: inst = 32'h24040000;
30'h00000141: inst = 32'h00042821;
30'h00000142: inst = 32'h00043821;
30'h00000143: inst = 32'h0c000023;
30'h00000144: inst = 32'h00000000;
30'h00000145: inst = 32'h3602f000;
30'h00000146: inst = 32'h8c420000;
30'h00000147: inst = 32'h00000000;
30'h00000148: inst = 32'h24030072;
30'h00000149: inst = 32'h0062182a;
30'h0000014a: inst = 32'h1460000e;
30'h0000014b: inst = 32'h00000000;
30'h0000014c: inst = 32'h24030061;
30'h0000014d: inst = 32'h10430018;
30'h0000014e: inst = 32'h00000000;
30'h0000014f: inst = 32'h24030064;
30'h00000150: inst = 32'h14430023;
30'h00000151: inst = 32'h00000000;
30'h00000152: inst = 32'h8fa70048;
30'h00000153: inst = 32'h00000000;
30'h00000154: inst = 32'h27a40050;
30'h00000155: inst = 32'h24050003;
30'h00000156: inst = 32'h24060000;
30'h00000157: inst = 32'h0800017a;
30'h00000158: inst = 32'h00000000;
30'h00000159: inst = 32'h24030073;
30'h0000015a: inst = 32'h10430012;
30'h0000015b: inst = 32'h00000000;
30'h0000015c: inst = 32'h24030077;
30'h0000015d: inst = 32'h14430016;
30'h0000015e: inst = 32'h00000000;
30'h0000015f: inst = 32'h8fa70048;
30'h00000160: inst = 32'h00000000;
30'h00000161: inst = 32'h27a40050;
30'h00000162: inst = 32'h24050000;
30'h00000163: inst = 32'h2406fffd;
30'h00000164: inst = 32'h0800017a;
30'h00000165: inst = 32'h00000000;
30'h00000166: inst = 32'h8fa70048;
30'h00000167: inst = 32'h00000000;
30'h00000168: inst = 32'h27a40050;
30'h00000169: inst = 32'h2405fffd;
30'h0000016a: inst = 32'h24060000;
30'h0000016b: inst = 32'h0800017a;
30'h0000016c: inst = 32'h00000000;
30'h0000016d: inst = 32'h8fa70048;
30'h0000016e: inst = 32'h00000000;
30'h0000016f: inst = 32'h27a40050;
30'h00000170: inst = 32'h24050000;
30'h00000171: inst = 32'h24060003;
30'h00000172: inst = 32'h0800017a;
30'h00000173: inst = 32'h00000000;
30'h00000174: inst = 32'hafa00044;
30'h00000175: inst = 32'h8fa70048;
30'h00000176: inst = 32'h00000000;
30'h00000177: inst = 32'h27a40050;
30'h00000178: inst = 32'h24050000;
30'h00000179: inst = 32'h00053021;
30'h0000017a: inst = 32'h0c000083;
30'h0000017b: inst = 32'h00000000;
30'h0000017c: inst = 32'h3c021bee;
30'h0000017d: inst = 32'h3c038000;
30'h0000017e: inst = 32'h24040070;
30'h0000017f: inst = 32'h3442f000;
30'h00000180: inst = 32'h34630020;
30'h00000181: inst = 32'hac440000;
30'h00000182: inst = 32'h8c620000;
30'h00000183: inst = 32'h00000000;
30'h00000184: inst = 32'h3c031800;
30'h00000185: inst = 32'hafa2003c;
30'h00000186: inst = 32'h8fa20040;
30'h00000187: inst = 32'h00000000;
30'h00000188: inst = 32'h34640004;
30'h00000189: inst = 32'hac820000;
30'h0000018a: inst = 32'h8fa20034;
30'h0000018b: inst = 32'h00000000;
30'h0000018c: inst = 32'h34630000;
30'h0000018d: inst = 32'hac620000;
30'h0000018e: inst = 32'h3c028000;
30'h0000018f: inst = 32'h34420020;
30'h00000190: inst = 32'h8c420000;
30'h00000191: inst = 32'h00000000;
30'h00000192: inst = 32'h8fa3003c;
30'h00000193: inst = 32'h00000000;
30'h00000194: inst = 32'h1043fff9;
30'h00000195: inst = 32'h00000000;
30'h00000196: inst = 32'h0800010e;
30'h00000197: inst = 32'h00000000;
30'h00000198: inst = 32'h00000190;
30'h00000199: inst = 32'h00000226;
default:      inst = 32'h00000000;
endcase
end
endmodule
